module N1(x,y,z);
   input y,z;
   output x;
   assign x = (y&z);
endmodule
